/* top.v */


module top (
    input wire btn,
    output wire led0,
);

    assign led0 = btn;

endmodule